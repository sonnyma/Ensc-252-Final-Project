LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
use work.definitions_package.all;

entity controlunit is
    port (
        clk, rst, hard_rst : in std_logic;
        inst : in std_logic_vector(2 downto 0);
		  toSeg : buffer arr8x5 := ("00000", "00000", "00000", "00000", "00000");
		  whenidle : out std_logic
    );
end controlunit;

architecture rtl of controlunit is

begin
	toSeg <= ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when ((rst = '1') or (hard_rst = '1')) else
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00010") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (inst = "001") and (rising_edge(clk))) else --message
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (inst = "010") and (rising_edge(clk))) else --snake to left
		("00011", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (inst = "011") and (rising_edge(clk))) else --snake to right
		("01000", "00000", "00000", "00000", "00000", "00000", "00000", "00110") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (inst = "100") and (rising_edge(clk))) else --fly
		("00000", "00000", "00000", "00000", "00000", "01101", "01110", "01110") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (inst = "101") and (rising_edge(clk))) else --error
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "01101", "01110", "01110") and (rising_edge(clk))) else --unerror
		("00000", "00000", "00000", "00000", "00000", "00000", "00010", "01111") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00010") and (rising_edge(clk))) else --half w
		("00000", "00000", "00000", "00000", "00000", "00010", "01111", "10000") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00010", "01111") and (rising_edge(clk))) else --w
		("00000", "00000", "00000", "00000", "00010", "01111", "10000", "10001") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00010", "01111", "10000") and (rising_edge(clk))) else --wh
		("00000", "00000", "00000", "00010", "01111", "10000", "10001", "10010") when (toSeg = ("00000", "00000", "00000", "00000", "00010", "01111", "10000", "10001") and (rising_edge(clk))) else --wha
		("00000", "00000", "00010", "01111", "10000", "10001", "10010", "00000") when (toSeg = ("00000", "00000", "00000", "00010", "01111", "10000", "10001", "10010") and (rising_edge(clk))) else --what
		("00000", "00010", "01111", "10000", "10001", "10010", "00000", "10011") when (toSeg = ("00000", "00000", "00010", "01111", "10000", "10001", "10010", "00000") and (rising_edge(clk))) else --what() 
		("00010", "01111", "10000", "10001", "10010", "00000", "10011", "10100") when (toSeg = ("00000", "00010", "01111", "10000", "10001", "10010", "00000", "10011") and (rising_edge(clk))) else --what d
		("01111", "10000", "10001", "10010", "00000", "10011", "10100", "10011") when (toSeg = ("00010", "01111", "10000", "10001", "10010", "00000", "10011", "10100") and (rising_edge(clk))) else --what di
		("10000", "10001", "10010", "00000", "10011", "10100", "10011", "00000") when (toSeg = ("01111", "10000", "10001", "10010", "00000", "10011", "10100", "10011") and (rising_edge(clk))) else --(half w)hat did
		("10001", "10010", "00000", "10011", "10100", "10011", "00000", "10010") when (toSeg = ("10000", "10001", "10010", "00000", "10011", "10100", "10011", "00000") and (rising_edge(clk))) else --hat did()
		("10010", "00000", "10011", "10100", "10011", "00000", "10010", "10000") when (toSeg = ("10001", "10010", "00000", "10011", "10100", "10011", "00000", "10010") and (rising_edge(clk))) else --at did t
		("00000", "10011", "10100", "10011", "00000", "10010", "10000", "01101") when (toSeg = ("10010", "00000", "10011", "10100", "10011", "00000", "10010", "10000") and (rising_edge(clk))) else --t did th
		("10011", "10100", "10011", "00000", "10010", "10000", "01101", "00000") when (toSeg = ("00000", "10011", "10100", "10011", "00000", "10010", "10000", "01101") and (rising_edge(clk))) else --()did the
		("10100", "10011", "00000", "10010", "10000", "01101", "00000", "10100") when (toSeg = ("10011", "10100", "10011", "00000", "10010", "10000", "01101", "00000") and (rising_edge(clk))) else --did the()
		("10011", "00000", "10010", "10000", "01101", "00000", "10100", "00000") when (toSeg = ("10100", "10011", "00000", "10010", "10000", "01101", "00000", "10100") and (rising_edge(clk))) else --id the 1
		("00000", "10010", "10000", "01101", "00000", "10100", "00000", "10101") when (toSeg = ("10011", "00000", "10010", "10000", "01101", "00000", "10100", "00000") and (rising_edge(clk))) else --d the 1()
		("10010", "10000", "01101", "00000", "10100", "00000", "10101", "10001") when (toSeg = ("00000", "10010", "10000", "01101", "00000", "10100", "00000", "10101") and (rising_edge(clk))) else --()the 1 s
		("10000", "01101", "00000", "10100", "00000", "10101", "10001", "10110") when (toSeg = ("10010", "10000", "01101", "00000", "10100", "00000", "10101", "10001") and (rising_edge(clk))) else --the 1 sa
		("01101", "00000", "10100", "00000", "10101", "10001", "10110", "00000") when (toSeg = ("10000", "01101", "00000", "10100", "00000", "10101", "10001", "10110") and (rising_edge(clk))) else --he 1 say
		("00000", "10100", "00000", "10101", "10001", "10110", "00000", "10010") when (toSeg = ("01101", "00000", "10100", "00000", "10101", "10001", "10110", "00000") and (rising_edge(clk))) else --e 1 say()
		("10100", "00000", "10101", "10001", "10110", "00000", "10010", "10111") when (toSeg = ("00000", "10100", "00000", "10101", "10001", "10110", "00000", "10010") and (rising_edge(clk))) else --()1 say t
		("00000", "10101", "10001", "10110", "00000", "10010", "10111", "00000") when (toSeg = ("10100", "00000", "10101", "10001", "10110", "00000", "10010", "10111") and (rising_edge(clk))) else --1 say to
		("10101", "10001", "10110", "00000", "10010", "10111", "00000", "10010") when (toSeg = ("00000", "10101", "10001", "10110", "00000", "10010", "10111", "00000") and (rising_edge(clk))) else --()say to()
		("10001", "10110", "00000", "10010", "10111", "00000", "10010", "10000") when (toSeg = ("10101", "10001", "10110", "00000", "10010", "10111", "00000", "10010") and (rising_edge(clk))) else --say to t
		("10110", "00000", "10010", "10111", "00000", "10010", "10000", "01101") when (toSeg = ("10001", "10110", "00000", "10010", "10111", "00000", "10010", "10000") and (rising_edge(clk))) else --ay to th
		("00000", "10010", "10111", "00000", "10010", "10000", "01101", "00000") when (toSeg = ("10110", "00000", "10010", "10111", "00000", "10010", "10000", "01101") and (rising_edge(clk))) else --y to the
		("10010", "10111", "00000", "10010", "10000", "01101", "00000", "10111") when (toSeg = ("00000", "10010", "10111", "00000", "10010", "10000", "01101", "00000") and (rising_edge(clk))) else --()to the()
		("10111", "00000", "10010", "10000", "01101", "00000", "10111", "11100") when (toSeg = ("10010", "10111", "00000", "10010", "10000", "01101", "00000", "10111") and (rising_edge(clk))) else --to the 0
		("00000", "10010", "10000", "01101", "00000", "10111", "11100", "00000") when (toSeg = ("10111", "00000", "10010", "10000", "01101", "00000", "10111", "11100") and (rising_edge(clk))) else --o the 0?
		("10010", "10000", "01101", "00000", "10111", "11100", "00000", "10101") when (toSeg = ("00000", "10010", "10000", "01101", "00000", "10111", "11100", "00000") and (rising_edge(clk))) else --()the 0?()
		("10000", "01101", "00000", "10111", "11100", "00000", "10101", "10010") when (toSeg = ("10010", "10000", "01101", "00000", "10111", "11100", "00000", "10101") and (rising_edge(clk))) else --the 0? S
		("01101", "00000", "10111", "11100", "00000", "10101", "10010", "10111") when (toSeg = ("10000", "01101", "00000", "10111", "11100", "00000", "10101", "10010") and (rising_edge(clk))) else --th 0? St
		("00000", "10111", "11100", "00000", "10101", "10010", "10111", "11000") when (toSeg = ("01101", "00000", "10111", "11100", "00000", "10101", "10010", "10111") and (rising_edge(clk))) else --h 0? Sto
		("10111", "11100", "00000", "10101", "10010", "10111", "11000", "00000") when (toSeg = ("00000", "10111", "11100", "00000", "10101", "10010", "10111", "11000") and (rising_edge(clk))) else --()0? Stop
		("11100", "00000", "10101", "10010", "10111", "11000", "00000", "11001") when (toSeg = ("10111", "11100", "00000", "10101", "10010", "10111", "11000", "00000") and (rising_edge(clk))) else --0? Stop()
		("00000", "10101", "10010", "10111", "11000", "00000", "11001", "10111") when (toSeg = ("11100", "00000", "10101", "10010", "10111", "11000", "00000", "11001") and (rising_edge(clk))) else --? Stop b
		("10101", "10010", "10111", "11000", "00000", "11001", "10111", "10111") when (toSeg = ("00000", "10101", "10010", "10111", "11000", "00000", "11001", "10111") and (rising_edge(clk))) else --()Stop bo
		("10010", "10111", "11000", "00000", "11001", "10111", "10111", "00010") when (toSeg = ("10101", "10010", "10111", "11000", "00000", "11001", "10111", "10111") and (rising_edge(clk))) else --Stop boo
		("10111", "11000", "00000", "11001", "10111", "10111", "00010", "01101") when (toSeg = ("10010", "10111", "11000", "00000", "11001", "10111", "10111", "00010") and (rising_edge(clk))) else --top bool
		("11000", "00000", "11001", "10111", "10111", "00010", "01101", "10001") when (toSeg = ("10111", "11000", "00000", "11001", "10111", "10111", "00010", "01101") and (rising_edge(clk))) else --op boole
		("00000", "11001", "10111", "10111", "00010", "01101", "10001", "11010") when (toSeg = ("11000", "00000", "11001", "10111", "10111", "00010", "01101", "10001") and (rising_edge(clk))) else --p boolea
		("11001", "10111", "10111", "00010", "01101", "10001", "11010", "00000") when (toSeg = ("00000", "11001", "10111", "10111", "00010", "01101", "10001", "11010") and (rising_edge(clk))) else --()boolean
		("10111", "10111", "00010", "01101", "10001", "11010", "00000", "11010") when (toSeg = ("11001", "10111", "10111", "00010", "01101", "10001", "11010", "00000") and (rising_edge(clk))) else --boolean()
		("10111", "00010", "01101", "10001", "11010", "00000", "11010", "11011") when (toSeg = ("10111", "10111", "00010", "01101", "10001", "11010", "00000", "11010") and (rising_edge(clk))) else --oolean (half m)
		("00010", "01101", "10001", "11010", "00000", "11010", "11011", "01101") when (toSeg = ("10111", "00010", "01101", "10001", "11010", "00000", "11010", "11011") and (rising_edge(clk))) else --olean m
		("01101", "10001", "11010", "00000", "11010", "11011", "01101", "00000") when (toSeg = ("00010", "01101", "10001", "11010", "00000", "11010", "11011", "01101") and (rising_edge(clk))) else --olean me
		("10001", "11010", "00000", "11010", "11011", "01101", "00000", "00000") when (toSeg = ("01101", "10001", "11010", "00000", "11010", "11011", "01101", "00000") and (rising_edge(clk))) else --lean me()
		("11010", "00000", "11010", "11011", "01101", "00000", "00000", "00000") when (toSeg = ("10001", "11010", "00000", "11010", "11011", "01101", "00000", "00000") and (rising_edge(clk))) else --ean me()()
		("00000", "11010", "11011", "01101", "00000", "00000", "00000", "00000") when (toSeg = ("11010", "00000", "11010", "11011", "01101", "00000", "00000", "00000") and (rising_edge(clk))) else --an me()()()
		("11010", "11011", "01101", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00000", "11010", "11011", "01101", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --n me()()()()
		("11011", "01101", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("11010", "11011", "01101", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --()me()()()()()
		("01101", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("11011", "01101", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --(half m)e()()()()()()
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("01101", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --e()()()()()()()
		("00000", "00000", "00000", "00000", "00000", "00000", "00001", "00101") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001") and (rising_edge(clk))) else --snake1 to left
		("00000", "00000", "00000", "00000", "00000", "00001", "00101", "00101") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00001", "00101") and (rising_edge(clk))) else --snake2
		("00000", "00000", "00000", "00000", "00001", "00101", "00101", "00010") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00001", "00101", "00101") and (rising_edge(clk))) else --snake3
		("00000", "00000", "00000", "00001", "00101", "00101", "00010", "00000") when (toSeg = ("00000", "00000", "00000", "00000", "00001", "00101", "00101", "00010") and (rising_edge(clk))) else --snake4
		("00000", "00000", "00001", "00101", "00101", "00010", "00000", "00000") when (toSeg = ("00000", "00000", "00000", "00001", "00101", "00101", "00010", "00000") and (rising_edge(clk))) else --snake5
		("00000", "00001", "00101", "00101", "00010", "00000", "00000", "00000") when (toSeg = ("00000", "00000", "00001", "00101", "00101", "00010", "00000", "00000") and (rising_edge(clk))) else --snake6
		("00001", "00101", "00101", "00010", "00000", "00000", "00000", "00000") when (toSeg = ("00000", "00001", "00101", "00101", "00010", "00000", "00000", "00000") and (rising_edge(clk))) else --snake7
		("00101", "00101", "00010", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00001", "00101", "00101", "00010", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake8
		("00101", "00010", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00101", "00101", "00010", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake9
		("00010", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00101", "00010", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake10
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00010", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake11
		("00101", "00011", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00011", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake1 to right
		("00101", "00101", "00011", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00101", "00011", "00000", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake2
		("00100", "00101", "00101", "00011", "00000", "00000", "00000", "00000") when (toSeg = ("00101", "00101", "00011", "00000", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake3
		("00000", "00100", "00101", "00101", "00011", "00000", "00000", "00000") when (toSeg = ("00100", "00101", "00101", "00011", "00000", "00000", "00000", "00000") and (rising_edge(clk))) else --snake4
		("00000", "00000", "00100", "00101", "00101", "00011", "00000", "00000") when (toSeg = ("00000", "00100", "00101", "00101", "00011", "00000", "00000", "00000") and (rising_edge(clk))) else --snake5
		("00000", "00000", "00000", "00100", "00101", "00101", "00011", "00000") when (toSeg = ("00000", "00000", "00100", "00101", "00101", "00011", "00000", "00000") and (rising_edge(clk))) else --snake6
		("00000", "00000", "00000", "00000", "00100", "00101", "00101", "00011") when (toSeg = ("00000", "00000", "00000", "00100", "00101", "00101", "00011", "00000") and (rising_edge(clk))) else --snake7
		("00000", "00000", "00000", "00000", "00000", "00100", "00101", "00101") when (toSeg = ("00000", "00000", "00000", "00000", "00100", "00101", "00101", "00011") and (rising_edge(clk))) else --snake8
		("00000", "00000", "00000", "00000", "00000", "00000", "00100", "00101") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00100", "00101", "00101") and (rising_edge(clk))) else --snake9
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00100") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00100", "00101") and (rising_edge(clk))) else --snake10
		("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000") when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00100") and (rising_edge(clk))) else --snake11
		("00111", "00000", "00000", "00000", "00000", "00000", "00000", "00111") when (toSeg = ("01000", "00000", "00000", "00000", "00000", "00000", "00000", "00110") and (rising_edge(clk))) else --fly1
		("00110", "00000", "00000", "00000", "00000", "00000", "00000", "01000") when (toSeg = ("00111", "00000", "00000", "00000", "00000", "00000", "00000", "00111") and (rising_edge(clk))) else --fly2
		("01100", "00000", "00000", "00000", "00000", "00000", "00000", "01001") when (toSeg = ("00110", "00000", "00000", "00000", "00000", "00000", "00000", "01000") and (rising_edge(clk))) else --fly3
		("01011", "00000", "00000", "00000", "00000", "00000", "00000", "00110") when (toSeg = ("01100", "00000", "00000", "00000", "00000", "00000", "00000", "01001") and (rising_edge(clk))) else --fly4
		("01010", "00000", "00000", "00000", "00000", "00000", "00000", "01010") when (toSeg = ("01011", "00000", "00000", "00000", "00000", "00000", "00000", "00110") and (rising_edge(clk))) else --fly5
		("00110", "00000", "00000", "00000", "00000", "00000", "00000", "01011") when (toSeg = ("01010", "00000", "00000", "00000", "00000", "00000", "00000", "01010") and (rising_edge(clk))) else --fly6
		("01001", "00000", "00000", "00000", "00000", "00000", "00000", "01100") when (toSeg = ("00110", "00000", "00000", "00000", "00000", "00000", "00000", "01011") and (rising_edge(clk))) else --fly7
		("00000", "01000", "00000", "00000", "00000", "00000", "00000", "00110") when (toSeg = ("01001", "00000", "00000", "00000", "00000", "00000", "00000", "01100") and (rising_edge(clk))) else --fly8
		("00000", "01000", "00000", "00000", "00000", "00000", "00110", "00000") when (toSeg = ("00000", "01000", "00000", "00000", "00000", "00000", "00000", "00110") and (rising_edge(clk))) else --fly9
		("00000", "00111", "00000", "00000", "00000", "00000", "00111", "00000") when (toSeg = ("00000", "01000", "00000", "00000", "00000", "00000", "00110", "00000") and (rising_edge(clk))) else --fly10
		("00000", "00110", "00000", "00000", "00000", "00000", "01000", "00000") when (toSeg = ("00000", "00111", "00000", "00000", "00000", "00000", "00111", "00000") and (rising_edge(clk))) else --fly11
		("00000", "01100", "00000", "00000", "00000", "00000", "01001", "00000") when (toSeg = ("00000", "00110", "00000", "00000", "00000", "00000", "01000", "00000") and (rising_edge(clk))) else --fly12
		("00000", "01011", "00000", "00000", "00000", "00000", "00110", "00000") when (toSeg = ("00000", "01100", "00000", "00000", "00000", "00000", "01001", "00000") and (rising_edge(clk))) else --fly13
		("00000", "01010", "00000", "00000", "00000", "00000", "01010", "00000") when (toSeg = ("00000", "01011", "00000", "00000", "00000", "00000", "00110", "00000") and (rising_edge(clk))) else --fly14
		("00000", "00110", "00000", "00000", "00000", "00000", "01011", "00000") when (toSeg = ("00000", "01010", "00000", "00000", "00000", "00000", "01010", "00000") and (rising_edge(clk))) else --fly15
		("00000", "01001", "00000", "00000", "00000", "00000", "01100", "00000") when (toSeg = ("00000", "00110", "00000", "00000", "00000", "00000", "01011", "00000") and (rising_edge(clk))) else --fly16
		("01000", "00000", "00000", "00000", "00000", "00000", "00110", "00000") when (toSeg = ("00000", "01001", "00000", "00000", "00000", "00000", "01100", "00000") and (rising_edge(clk))) else --fly17
		("01000", "00000", "00000", "00000", "00000", "00000", "00000", "00110") when (toSeg = ("01000", "00000", "00000", "00000", "00000", "00000", "00110", "00000") and (rising_edge(clk))); --fly18

	--to check when a program finishes (makes 1 when at the end of program, else 0)
	whenidle <= '1' when (toSeg = ("01101", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (falling_edge(clk))) else
		         '1' when (toSeg = ("00000", "01001", "00000", "00000", "00000", "00000", "01100", "00000") and (falling_edge(clk))) else
					'1' when (toSeg = ("00000", "00000", "00000", "00000", "00000", "00000", "00000", "00100") and (falling_edge(clk))) else
					'1' when (toSeg = ("00010", "00000", "00000", "00000", "00000", "00000", "00000", "00000") and (falling_edge(clk))) else
					'0' when falling_edge(clk);
end architecture;