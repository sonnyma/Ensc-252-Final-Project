library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity snake is
    port (
        clk : in std_logic;
        rst : in std_logic;
    );
end snake;

architecture rtl of snake is

begin

end architecture;