library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity message is
    port (
        clk : in std_logic;
        rst : in std_logic);
end message;

architecture rtl of message is

begin

end architecture;