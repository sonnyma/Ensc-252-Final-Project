library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fly is
    port (
        clk : in std_logic;
        rst : in std_logic;
    );
end fly;

architecture rtl of fly is

begin

    
end architecture;